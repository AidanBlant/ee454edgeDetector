
module threshold #(parameter WIDTH, parameter DEPTH)(
	input threshold,
	input [WIDTH*DEPTH:0] inputImage,
	output outputImage
);



initial
begin

	
end

endmodule